Gena
True
228
